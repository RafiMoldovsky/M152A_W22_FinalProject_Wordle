module word_db (input [24:0] word, output wire in_db);

//Bloom filter storing 1000 words in 4096 bits with 4 hash functions
localparam [11:0] hash_params [0:3] [0:4] = {
{12'h0dcb, 12'h05bc, 12'h0adf, 12'h0dd2, 12'h021c},
{12'h0869, 12'h037a, 12'h08b5, 12'h0566, 12'h0a69},
{12'h0613, 12'h0641, 12'h0fc8, 12'h0d28, 12'h04cf},
{12'h0c66, 12'h0602, 12'h025c, 12'h0387, 12'h0a6f}
};

(* ramstyle = "block" *) localparam bloom_filter [0:4095] = {
64'b111011111100100010010101101100110101101100110100110111110100110,
64'b100011101111101001111100011011110101111001100101101011111101111,
64'b110111101101100111111111100011110011111001111111010111110111110,
64'b011111101110110110000111011011111100000101101111111001100101100,
64'b111011010110110100110111100000011100111111111111110010101011001,
64'b111111000001011011011110001110111111101101100111000011011000001,
64'b000111000000011101111110001110110101111101110101101000001101000,
64'b111001101011010011111010111000110000110111111100111111001101111,
64'b011011011000011111101101000101101111110111110100011111111110110,
64'b100111111001101101101010110111111001001110010110110101011011110,
64'b011101001100001101011111011011010100011110101111101000010001111,
64'b011111111111010111111001010111011111101101101011010010101111101,
64'b101011000111001111011101100110110110101101110111100011001111000,
64'b111111011111001011100111111111011001011111100100111011000101010,
64'b101101100101010101110111111110011111100000010110010111011010111,
64'b010011011110100101010100111110011010001000111110110100110101011,
64'b101110110111110101010111100111111000011101111110111011011101111,
64'b111000111101101001011100101101100101111100100001011111110000111,
64'b111111111010110111111110000101111101101111101010111111011111101,
64'b110001011111110111110001011100011001010001010011101111011110101,
64'b110110011010111111010110100001100010110011111010111111011011001,
64'b010110111010011011001011011101010111011101000000011101111101111,
64'b110010110110011111101111111110111111101110111111100011111110111,
64'b000110110001100111001000100001111011110100110110010010011000111,
64'b100101101011000011010111010010110111110111000110111111100111011,
64'b110111010110101101110111010110000111011011011001101111111011100,
64'b110111100001011011111110010101111111000010001101111101100101011,
64'b110100110000111111010010111111100111111100111111100011110110101,
64'b101111110001110111111011011010011110011110111111101101111101010,
64'b111101000110010111110111110011011101101111010111110110111011010,
64'b101111111010010011111111001101110011011001010110100100111011001,
64'b111101000001101011110110010101011111010011010001010110111100010,
64'b101011000100101110010101011011111011111001110101000001010110101,
64'b010100110100011110111010011111001010011111101110111010011001011,
64'b100010001010110011011001111110111111111111010101000111001011110,
64'b010011011100011101001101100111101111111010111110111010111011110,
64'b011110101101011111111001011011101111011101110010101111111101011,
64'b011101000001110111011110111100110111101010001101010111001010111,
64'b110101100111111101101101111011100111100101000010110011110010001,
64'b011001111011001011111111001100111111101111011111101100100010110,
64'b010101000111010001100000101001011010111101011100110101101110011,
64'b001011111101001111101001001100101111110111111001010111101010001,
64'b111110110000110111110110011011100010001111011100110111001010110,
64'b111101011101011010011001011101000101010100110101110011010010000,
64'b100010111111111111011111000011100111110110101011110010100011010,
64'b111011001111100010001111111101001111001101001110010111010011000,
64'b111011011111101010101101110001000110101000001111111111011110100,
64'b101011001010101100100101101100011101111111010111110111010011111,
64'b010111111000110001100111001111111101101001010111111001101101011,
64'b100110010001110111111111110010001111011110111101011100011101011,
64'b111110011011110111011111110010111010110010111110000011101111110,
64'b011011110000111000010111110001111101010100000101011010101100011,
64'b101110111001010011101111001111011011001100111101110010101011110,
64'b011100011011100111000110011110100011100010110111010011100110111,
64'b110011110110101101111110110110111101011110001011001011101101010,
64'b110100100101101101110010011001110000101001110110110101101010011,
64'b100100000010101111000011010111110111100011110111110110011001010,
64'b110101101011011011010111111010101101101111111100010100000001010,
64'b111111001100001001111110110001001101111110100001000100110010001,
64'b111111111111101001111010001010010101111101001111111011100011000,
64'b110011010111111110011100110011111110101101011110110110111111011,
64'b111010000111111001011100110100100110111111011111010100100110101,
64'b001110011010111011101010000111010110110001101011011010101110111,
64'b111101010001111111111110110110101111010001101111100101110110100
};

wire [11:0] hash_table [0:4];

wire [11:0] hash;

reg [0:3] in_db_i;

reg [1:0] i;

genvar j;
generate
for (j = 0; j < 5; j = j + 1) begin : which_letter
assign hash_table[j] = hash_params[i][j] * word[5*j + 4:5*j];
end
endgenerate
assign hash = hash_table[0] + hash_table[1] + hash_table[2] + hash_table[3] + hash_table[4];

always @(posedge clk or posedge rst) begin
    if (rst) begin
        i <= 0;
        in_db_i <= 4'b0;
    else begin
        i <= i+1;
    end
end
        
assign in_db_i[i] = bloom_filter[hash[i]];

assign in_db = &in_db_i;

endmodule
