module target_word(input [6:0] index, output [24:0] word);

localparam [24:0] wordlist [0:99] = {
25'b1001110110001000000001010, //tweak
25'b0000110001001000000001010, //break
25'b0100101110010100010010001, //joker
25'b0101100000000110101100100, //ladle
25'b0011001000000000110110011, //giant
25'b0010001101100111000111000, //entry
25'b1001001110010111010100100, //solve
25'b0010001011101000001100100, //elude
25'b1001010110001000000010011, //sweat
25'b0011100000100011000111000, //harry
25'b0001100100100110111010111, //detox
25'b0101101110101100101111000, //lowly
25'b0010110001011100110100011, //frond
25'b0001010001001000010001010, //creek
25'b1001000111010001000101010, //shirk
25'b0001000000011110010010001, //caper
25'b0011101110000010000111000, //hobby
25'b0000101011011100111001100, //bloom
25'b0101101110101001001011000, //lousy
25'b0110001110101000101110011, //moult
25'b0011101000011010011000100, //hinge
25'b0001101000100111001111000, //ditty
25'b0011010100000001010100000, //guava
25'b1011001110100011000111000, //worry
25'b1001100000011110010010001, //taper
25'b0010101011010000110110011, //flint
25'b0010000001011100110111000, //ebony
25'b0101101110000000110011000, //loamy
25'b0110101110100011001100111, //north
25'b0001100100000010100010011, //debit
25'b0010101011101001001000111, //flush
25'b0110100100101010010010001, //never
25'b0001100100000011010010011, //debut
25'b0110001000000101000101110, //micro
25'b0000010001001000110100000, //arena
25'b0110010100100100011111000, //mushy
25'b0111101011000001001100100, //plate
25'b0001010001001001001010011, //crest
25'b0110101000001000001000100, //niece
25'b1001000111000001011001011, //shawl
25'b0001010001011101011001101, //crown
25'b1001000111010000110100100, //shine
25'b0000100000011010000001011, //banal
25'b0000000110000001001100100, //agate
25'b0111010100100110010010001, //outer
25'b0001110001010001010100100, //drive
25'b1001010100100010010010001, //surer
25'b0011000000101000011000100, //gauge
25'b0010101000000101010010010, //ficus
25'b1001110001010000001000100, //trice
25'b0110001110100101001011000, //mossy
25'b0110101110010001001011000, //noisy
25'b0000101011000000110101010, //blank
25'b1001000000010111010101110, //salvo
25'b0001110110000001000100101, //dwarf
25'b0111100000010111001011000, //palsy
25'b0011001110000110101111000, //godly
25'b0010100100011000110000100, //femme
25'b1001000111010000010110011, //shift
25'b0010101011011100111010001, //floor
25'b0010101000001011001111000, //fifty
25'b1000010100000000001001010, //quack
25'b1001010011000001001000111, //stash
25'b0001010001001000000001010, //creak
25'b1010001101001010100010011, //unfit
25'b0110000100010110010000100, //melee
25'b0101111000011010001000111, //lynch
25'b0110000000011010100000000, //mania
25'b1001000111011100111010011, //shoot
25'b1010100000010111010000100, //value
25'b1001000100101010010001101, //seven
25'b1001100000010100010001101, //taken
25'b1000100100000011010010011, //rebut
25'b0111100000100010010010001, //parer
25'b0011001011011100000100100, //globe
25'b1001100111110000110000100, //thyme
25'b0001101000101010010010001, //diver
25'b1001001011101001000101111, //slurp
25'b0001110001000000100001101, //drain
25'b1001110110010001011110011, //twixt
25'b0110010100100010000001011, //mural
25'b1001100000101100110111000, //tawny
25'b1001000010000000101101111, //scalp
25'b1001001111100010010000100, //spree
25'b1011001110100010101100011, //world
25'b0000000111001000000000011, //ahead
25'b1011010001101000110100110, //wrung
25'b0001010001001000110000100, //creme
25'b1011001000100100010010001, //wiser
25'b0001000000100010011001110, //cargo
25'b0111110100100011001000100, //purse
25'b1001000111001000010010011, //sheet
25'b0111010101010000110100100, //ovine
25'b0101101000010110000000010, //lilac
25'b0000001100010001001111000, //amity
25'b0111100111011100110100100, //phone
25'b0001001110011010100000010, //conic
25'b1001000111110000101111000, //shyly
25'b0101100100000000010111000, //leafy
25'b0110001110101100010010001 //mower
};

assign word = wordlist[index];

endmodule
