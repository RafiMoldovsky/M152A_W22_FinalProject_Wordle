`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:30:38 03/19/2013 
// Design Name: 
// Module Name:    vga648'h480 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vga640x480(
	input wire dclk,			//pixel clock: 25MHz
	input wire clr,			//asynchronous reset
	output wire hsync,		//horizontal sync out
	output wire vsync,		//vertical sync out
	output reg [2:0] red,	//red vga output
	output reg [2:0] green, //green vga output
	output reg [1:0] blue	//blue vga output
	);

// video structure constants
parameter hpixels = 800;// horizontal pixels per line
parameter vlines = 521; // vertical lines per frame
parameter hpulse = 96; 	// hsync pulse length
parameter vpulse = 2; 	// vsync pulse length
parameter hbp = 144; 	// end of horizontal back porch
parameter hfp = 784; 	// beginning of horizontal front porch
parameter vbp = 31; 		// end of vertical back porch
parameter vfp = 511; 	// beginning of vertical front porch
// active horizontal video is therefore: 784 - 144 = 640
// active vertical video is therefore: 511 - 31 = 480

// registers for storing the horizontal & vertical counters
reg [9:0] hc;
reg [9:0] vc;

// alphabet bitmaps
// ARTWORK
localparam ALPHABET [0:25][0:7][0:7] = {
	 { 8'h0C, 8'h1E, 8'h33, 8'h33, 8'h3F, 8'h33, 8'h33, 8'h00},   // U+0041 (A)
    { 8'h3F, 8'h66, 8'h66, 8'h3E, 8'h66, 8'h66, 8'h3F, 8'h00},   // U+0042 (B)
    { 8'h3C, 8'h66, 8'h03, 8'h03, 8'h03, 8'h66, 8'h3C, 8'h00},   // U+0043 (C)
    { 8'h1F, 8'h36, 8'h66, 8'h66, 8'h66, 8'h36, 8'h1F, 8'h00},   // U+0044 (D)
    { 8'h7F, 8'h46, 8'h16, 8'h1E, 8'h16, 8'h46, 8'h7F, 8'h00},   // U+0045 (E)
    { 8'h7F, 8'h46, 8'h16, 8'h1E, 8'h16, 8'h06, 8'h0F, 8'h00},   // U+0046 (F)
    { 8'h3C, 8'h66, 8'h03, 8'h03, 8'h73, 8'h66, 8'h7C, 8'h00},   // U+0047 (G)
    { 8'h33, 8'h33, 8'h33, 8'h3F, 8'h33, 8'h33, 8'h33, 8'h00},   // U+0048 (H)
    { 8'h1E, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h1E, 8'h00},   // U+0049 (I)
    { 8'h78, 8'h30, 8'h30, 8'h30, 8'h33, 8'h33, 8'h1E, 8'h00},   // U+004A (J)
    { 8'h67, 8'h66, 8'h36, 8'h1E, 8'h36, 8'h66, 8'h67, 8'h00},   // U+004B (K)
    { 8'h0F, 8'h06, 8'h06, 8'h06, 8'h46, 8'h66, 8'h7F, 8'h00},   // U+004C (L)
    { 8'h63, 8'h77, 8'h7F, 8'h7F, 8'h6B, 8'h63, 8'h63, 8'h00},   // U+004D (M)
    { 8'h63, 8'h67, 8'h6F, 8'h7B, 8'h73, 8'h63, 8'h63, 8'h00},   // U+004E (N)
    { 8'h1C, 8'h36, 8'h63, 8'h63, 8'h63, 8'h36, 8'h1C, 8'h00},   // U+004F (O)
    { 8'h3F, 8'h66, 8'h66, 8'h3E, 8'h06, 8'h06, 8'h0F, 8'h00},   // U+0050 (P)
    { 8'h1E, 8'h33, 8'h33, 8'h33, 8'h3B, 8'h1E, 8'h38, 8'h00},   // U+0051 (Q)
    { 8'h3F, 8'h66, 8'h66, 8'h3E, 8'h36, 8'h66, 8'h67, 8'h00},   // U+0052 (R)
    { 8'h1E, 8'h33, 8'h07, 8'h0E, 8'h38, 8'h33, 8'h1E, 8'h00},   // U+0053 (S)
    { 8'h3F, 8'h2D, 8'h0C, 8'h0C, 8'h0C, 8'h0C, 8'h1E, 8'h00},   // U+0054 (T)
    { 8'h33, 8'h33, 8'h33, 8'h33, 8'h33, 8'h33, 8'h3F, 8'h00},   // U+0055 (U)
    { 8'h33, 8'h33, 8'h33, 8'h33, 8'h33, 8'h1E, 8'h0C, 8'h00},   // U+0056 (V)
    { 8'h63, 8'h63, 8'h63, 8'h6B, 8'h7F, 8'h77, 8'h63, 8'h00},   // U+0057 (W)
    { 8'h63, 8'h63, 8'h36, 8'h1C, 8'h1C, 8'h36, 8'h63, 8'h00},   // U+0058 (X)
    { 8'h33, 8'h33, 8'h33, 8'h1E, 8'h0C, 8'h0C, 8'h1E, 8'h00},   // U+0059 (Y)
    { 8'h7F, 8'h63, 8'h31, 8'h18, 8'h4C, 8'h66, 8'h7F, 8'h00}   // U+005A (Z)
};

 reg [31:0] ctr;
 always @(posedge dclk) begin
 ctr <= ctr + 1;
end

wire in_db;

word_db Word_db(.word(ctr), .in_db(in_db));

// Horizontal & vertical counters --
// this is how we keep track of where we are on the screen.
// ------------------------
// Sequential "always block", which is a block that is
// only triggered on signal transitions or "edges".
// posedge = rising edge  &  negedge = falling edge
// Assignment statements can only be used on type "reg" and need to be of the "non-blocking" type: <=
always @(posedge dclk or posedge clr)
begin
	// reset condition
	if (clr == 1)
	begin
		hc <= 0;
		vc <= 0;
	end
	else
	begin
		// keep counting until the end of the line
		if (hc < hpixels - 1)
			hc <= hc + 1;
		else
		// When we hit the end of the line, reset the horizontal
		// counter and increment the vertical counter.
		// If vertical counter is at the end of the frame, then
		// reset that one too.
		begin
			hc <= 0;
			if (vc < vlines - 1)
				vc <= vc + 1;
			else
				vc <= 0;
		end
		
	end
end

wire box_i;
assign box_i = (vc - vbp) / 80;

wire box_j;
assign box_j = (hc - hbp - 120) / 80;

wire [2:0] ltr_x;
assign ltr_x = ((vc - vbp + 72) % 80) / 8;
wire [2:0] ltr_y;
assign ltr_y = ((hc - hbp + 32) % 80) / 8;

wire v_in_box;
assign v_in_box = ((vc - vbp + 72) % 80) < 64;

wire h_in_box;
assign h_in_box = ((hc - hbp + 32) % 80) < 64;


// generate sync pulses (active low)
// ----------------
// "assign" statements are a quick way to
// give values to variables of type: wire
assign hsync = (hc < hpulse) ? 0:1;
assign vsync = (vc < vpulse) ? 0:1;

always @(*) begin
// first check if we're within vertical active video range
	if (vc >= vbp && vc < vfp)
	begin
		// main display area
		if (hc >= (hbp) && hc < (hbp+640))
		begin
			// main game area
			if (hc >= (hbp+120) && hc < (hbp+520)) begin
				if (h_in_box && v_in_box) begin
					if (ALPHABET[box_i + box_j][ltr_x][ltr_y]) begin
						red = 0;
						green = 0;
						blue = 0;
					end else begin
						red = 3'b111;
						green = 3'b111;
						blue = 2'b11;
					end
				end else begin
					red = 0;
					green = 0;
					blue = 0;
				end
			end
			// Ukraine flag
			else if (vc >= (vbp + 240)) begin
				red = 3'b111;
				green = 3'b111;
				blue = 0;
			end else begin
				red = 0;
				green = 0;
				blue = 2'b11;
			end
		end
		// we're outside active horizontal range so display black
		else
		begin
			red = 0;
			green = 0;
			blue = 0;
		end
	end
	// we're outside active vertical range so display black
	else
	begin
		red = 0;
		green = 0;
		blue = 0;
	end
end

endmodule



//Bloom filter storing 5757 words in 32768 bits with 4 hash functions
localparam [14:0] hash_params [0:3] [0:4] = {
{15'h3aba, 15'h5b55, 15'h66ba, 15'h4f75, 15'h1093},
{15'h76f4, 15'h3092, 15'h5d56, 15'h0cb7, 15'h263b},
{15'h0d13, 15'h128d, 15'h56d3, 15'h0c5a, 15'h374f},
{15'h3643, 15'h36ac, 15'h5a38, 15'h1ae7, 15'h4334},
};
localparam [32767:0] bloom_filter = {
128'b0011111001010110101110011011111011010101111110101101011001010110111101111001100001011110111000100100011001010100110010100010001,
128'b1010111101101100101100111101111011101111010011011101110100000110011011001010011001101000000000000000100001010011010100100111000,
128'b1001101100110111010101101101001111001000010101101001001011000110101010110101010000101110000010111010000001001111101100111011101,
128'b1000111010101000111101101000111000010011100110011000111010111010111011101000111010111111000000110110010110111011000111011001100,
128'b0101011001011001100011110111000011111111100111110011110011100011001111001111001111001111011101100111001101110100010001101101011,
128'b0011000000011101111000011011101100110100000011111011011100001001001110011001111110101111100101100010110011110010111100111110001,
128'b0111101011100011110010001001100100001111101010111001110100101010010101111011010110100101110111100110010100111010000011001000001,
128'b1100000110100010110011101000000110111110101101001110001101100100010001001101111101110111101110011001100000100010001000000101011,
128'b0100110000110111101001000110001111001100000011111001111010110001111111011010111111010101101110010100101000101111000001001100001,
128'b0010010110110101101001010001000001100100001101001011101100010000000100000101001101100100100011111101110100000110001101110111100,
128'b1010001000010011010110000110000001011101000101110101100111111100101000111101101001110111011111110010111010011000111111101111110,
128'b1000110101111010000100110111011100000000110100011000011111111010110011010010010011000101011001110010101100100011001010000011110,
128'b1010001111010001111111010100000111011000011000101000010100001100111000100101100100111111010000001101111010110001101100010010101,
128'b0011111101110001100110000000001010100110101110101001001111100000101001111001000111001010011111110100101100011011111011110101010,
128'b1110010111001101110101011101100111110101011010101010110011110111101100100101111111110110000001100000010110000100110110011000110,
128'b0010100000110101010001110101010100001000000110101101010000111011111111001101011010101101011101100001111000011000111110000110111,
128'b0111110100001011111010010111010010001110011100010010011101110100100110110111001001011011001111010000010011101101001000010100110,
128'b1000001101011000101000010110011001001000000100001000110110011011001000010000010110000000001010011110101011110011011110110100010,
128'b1000010000110011101110000011111111111111011011010010001000100111000011110110101010101110101000001001111110000000010101111100101,
128'b0001001100001010000010110000000111100111111000010111111010110010110001110111110110111000010111100101010001111100010100111100111,
128'b1101101010010110100000000110110001000000101110010110110001101011000101000101011101110011010010100111000011111010110000000010001,
128'b1011100111101111101010110000011101110000001010001101111010000101100100010001111101100001011110001000111110000101111101101111010,
128'b1011011011001110101110010000101000000001100000001011010011010111110000011110101000010001000000111110010001101101110001101010101,
128'b1010010110010001100101101100011010110111011001101000101011000001010100001010111000111111001001100100011101100110001100001011011,
128'b1001000011110000011000110110001110010011010100000111110001000110111110010011000001010010111010100111000111010001010000001110111,
128'b1101011011110111100001010011000110011000100100010110001101000101010110010101110111010110110010000101000110000111010100111000001,
128'b0110110010110111011111011101100010001010100000000000000001111110111101110111000101111101101100100010111111010100010001001001011,
128'b0000011011101111101001011101010001111000001000111011011111100101001000010100110010110010101101011010101000001001111100111011001,
128'b0101000001100100110100001110100110100100101010111111001010010010000011100101010100010111001111001011100100001011111101011010111,
128'b1011000100111111101010001100100001011011000111011111100011111001001111000111001000000011001010011010111101100110001100111001100,
128'b0111111011011011101000010101010010000101011001110101011100001001100100010100101010101100010011111010011101010100010010010100011,
128'b0100110010000100110011101000001100110111010001100011101100000001001000101011110010000110000001110001010000111001000111110000101,
128'b0000000001010110101000000101100010010101101111010000100011000100110001011101011101010110011011101000110011110100010100001101010,
128'b0001001000101000000111011110011100110001010010011101011110001111011010101001011001110110010011011011011001110010001111000100001,
128'b0101110011010100010101110010110101000111111000010111001000110010111100110100010100110100010100001111011011100101110111000110010,
128'b1111001101101101011101001111011010110101110111001100010010101100000101011000011000000110110111111011011101011111011010110000011,
128'b0001111110000111010001001100111111000000010100010010110010010111111100011101110100010110001110011100011100010011110111000100000,
128'b0101011110110010100110100010010110000110101011101101101011010001011001010110110001110100110101110101100111001101101011110011110,
128'b0010010111110111110001001100100010110100010001010010101001100001011110010011001011100000000111000000011001010011010100001011101,
128'b1101101010110110110000100111110100100111011100010101010001111101111111001010111100000011100101011111110000110100100001000111110,
128'b1111110001001100111101111111010000001000110010110110100100000101011010011110011001001101001010010110000110100000101111111101100,
128'b1110010001111100101110100010100001010100000010010001000101101110100111010111011001111011011110001000110101100111010001011111111,
128'b0011010110111010001001110111110111000001011011111111000000010100101001111100110011001101111011000000001100010101111101111111100,
128'b1001010111111101010100000101110011111011100100010000111111000100100110100011011110010010011000000010111001101110000111011000110,
128'b1011111011001101100111101001010000011000111110101010110010011100100000000101010010110010101110110100001000010101111000111010001,
128'b0001100000111100011010111010010001010000111100101101010100001110010001011001110111111100001000000101010111101100110111011101001,
128'b1100111010101110111101010000111111101001011000100101111011010101001011000110100101001111111110000010010111010111111010010110111,
128'b0011100110111001000011101000101110000111101110110011000010100100110101100101111110010110000110000010100010111011000010111100110,
128'b0010100101100110110001011011000100010101001100010101111101010001010001010000100010110110100111001111001110100101000111010001010,
128'b0110111111010000000110110001000010001011000001000001011101101100110110011011000100100000100011111110011101110100111010001111000,
128'b1100111010010010001011000011110001000101011000000100011101110100100001010001000111011111111011011010001011000100000001001100111,
128'b1111011111001110111011100111110111011111001110110101000101101011011110001111110100111000110011000010000111011111101000011000111,
128'b0010111001110111111001101011010011000011000101000010011111001110111101101010110010000100011010111011101000111011101011000001010,
128'b0101101110110001000011011011101110100111100111001001110101011100101001110111001010010111111100011011100010111001010011101100011,
128'b1000011001111100110111001111100010110010001011101111000100110101101100010001111000000001001010110110100000111011000001010110101,
128'b0110010101110011000010011000101100111110010110010101110100100011000001101000010111110001001001111011100000100100010110010101101,
128'b1001001111111000101100100101011001111100110111100101010000100100111011101100011011111001101110101011011100010110011001100110010,
128'b0000101011111111000100110100101111010110010101110011010010001110000011001101111011110001100010111101011100001111111100000110110,
128'b1000101010111010111000011100010010100110010110000001001101100011101101111111000011001100001011101101100000010101110101000011100,
128'b0110101000001110100111101100011110011011000101011110010000001011001001000101101000100001111110011011001111011111001000111010111,
128'b0110001001101110001001111011011111001000110101011101100111101101111101101111111000111110010100111101001101100100100010000110010,
128'b0011010000000011011011110010001011101111000010101000001000010100011111100101001010110110011011010010010111100111110100010111001,
128'b1010111000001100100101101001011101010011100101101000100000100101101111010011001000000110011101000011010010011101011000110011110,
128'b1101110111010110111100111011001000101110110100011110010101100011110101110110110110000111001111111011001101110111101111111111101,
128'b0010111001010000100011100001001101100011110100111011111100101111001010110010001001011010010001001010100000010100101101001010001,
128'b1011010001110101011001011101010000010001000011100110101001000110011011111001111010001101001100011100011011010101111101000000001,
128'b1001100001110110100100011101010101100000000001110010010010001000001000100110101001001000100000001100000000101101010100110000111,
128'b0011100001101100010111100011011000100100001111100010000101110101101110001110101110100100000011101101010001100101111010011001000,
128'b0000111101001011111110000100001001010001101000001010010100011010000011111101000100111100010101100000011010010101100110111101000,
128'b0000111111000000010001100001000111010111100001010001001010110110111010101111000111111011010111100101001110001010011101101101111,
128'b1111010001110101110110010000011001110001100001011111001110100100010011101111000001011100010100101000100000010111001001100011011,
128'b0100110000100110101001011110000001110111010110110011001001000111010101001100000100000110100101111000110010110100010000001110010,
128'b0110000100011110110111110101101100000111011100000000010110111101111000001011011001011111110010001110011001110100011011001001010,
128'b1000110111001101101101010100000011110100100001100101101111011011101110101110010101100000001111001000110001001000110101001000111,
128'b1100100110010011000010111000010000100101110101110110011101111100100011001101000000011111100010000011011001011011011100111001010,
128'b1100100001100100101100110111001011010111111011010101000110110010101100010011100011101010101101000001110111000000000101000101001,
128'b1011110100010001111101010100101011100101110011100010101011010000010110001011001111000011000001011001001101110110101001110000110,
128'b0001000111001100000100001000100100110010100011010001010001101000000110111100110000011010100000110100011111111100000101000001010,
128'b1001010100001011101111010010111000000001010111011010011110110110011010011001000100000001010110001011110101101100100100011001101,
128'b0000000000000100011011010001100000001000101010110101001010000100111101001011010111011101010111101100010001101011101001100001110,
128'b0011111110011010111110100111001011111001010001011101111000001111101001000111110000110101100010000011110110111111010000100001111,
128'b0001101111001110110011101001010111100100110000001010110001101111101111110010111011001100111000110011010100111100101110101011011,
128'b0110100110010010001011111111100000011001100111001010011101000111100110000011111011010010011101101001100001101010010000001110101,
128'b1111011001110010010011011000101101001000110010001011100000010110001111000001010111001100000101000111011110100011111110000110000,
128'b0110100101100101001110110110001000010011010100110010101110011111000011110011010110110110111100001111010110011010001011011110110,
128'b0111011111100101100001010111000101001000001110110111010000011110000110000000110111011100000100101111100110010001001001100110101,
128'b0110101110010000101100001111100100100011110010011111011011011110101100111011011110010010000111101010111111010100110110110001001,
128'b1000001010001001001111000100011000001001111011010110010111110110110101110101100101110101100110001100110111011111010010101011010,
128'b0011000100111001111100100100111011001111100001010100111000101001011000001111011111110111000010101100010111000101110111110111011,
128'b1111111110101011100101010101001110010010010001001101001101100010011111101100111011010000101010110011111101010001110100001011010,
128'b0001101100010000101101101010010010110001101010010110100101111011111100111111110000111110010101100110001011111010101010001001010,
128'b0100001000101101110000011010001100101110100010010010000001010001000000000111110100111110111000111001111110011101100101000100101,
128'b1110100111011011111110111111110000100011111110100110100001110111010110010000000100101111011000000010011101010100110101111101101,
128'b0110011011110100011100000111011011111000001001000101011101101001001101101001111000110011110110010110010110110110101000010010000,
128'b1110111011011100100111000011011111111111100100100010110000101111111111111110000101101001110111100100111110111101011011111011010,
128'b0011110000000011000100011101101100111010110010011000101001101101000111101001110100011111011011101000000011010100000111101100011,
128'b1110100110100000001101110011000011101110010110100001001001110100011010101100100000000011110100000100101011001011000000110001011,
128'b0001011000101101010100010001011000111111010101001010000000111100010000110100010010100100011111110010111100110110011111010000100,
128'b1110111010011000111101110000011110101011111010000011110100000010101011110001000011111000110110011110100100110101111010100000001,
128'b0000000100110110011101000111110011001111110100110010111101010101111110100000101001010011000100001011100110000001110101111101011,
128'b1000000100011111100100011001001001011100011010111110001010010100110100001110111110010000001000001011000000111011110001011101111,
128'b0010011101110101000011000101010111110100100011000100111111011011110001011111110101111001001000110111011111001000011010111110001,
128'b1000001010010011000000110100000101111110101001000101111001111010101101110001000110001011000001110001111010011101010111001111110,
128'b1100110110010001100111010111101101100111101111010011000101011110001000111110101010110001110100011110110110010101101100101011100,
128'b1111011001011100000000010001000110011101000111110100000000010101010101100001011100111011100110110011011100001100110110000101100,
128'b0011011011000100001010110100001010001111011001011101101000100111001011010001001100001001011011010010110100000001001010100100011,
128'b1111001001100011011101101101001110010001001011010110100110111100110010101011111100001110101110001000010110111011011000110010110,
128'b0111011000111001010101111110011110010111100110111110111000010111101100000110010001100010100001001100000001010101110110111001111,
128'b0111111100100110111110010001011101101110001111010111111010010001010011011011100110000111010010001001000001010111110101011100011,
128'b0011111111110010000111010001000011100010000010011110101110010010110001101000101011110000000111011101100111111011101100110101010,
128'b1010000111110111001010000100000010100001001100111110010011000110010111110101000101001000001011110111010011001000101110000110001,
128'b0011010111001101011010000001101101000101001101010001111001101111010100001001110001111001001001111110010010100100011110110111101,
128'b1110101100100000011110101101001101110011010110111000010000111101111011011100011111010001111001101000010001000010010111111011000,
128'b0010110111101100000111000000000100100011110101100010011001001100001100101101111110111101011011111111000010110011011111111111001,
128'b0011001001001111010100110111001100001111010101010010101100111100010011000101100000111000011010010101100011011100101010111100100,
128'b0111011111100000011010001111001111010100011000100110000011001011101011101000111101101110110100001011011100101000110011010110011,
128'b1011010101011111110110001111011110000001101110010101010101101100001110011000111111100000101010011011010111101100011111000010001,
128'b1101100010010101111001010001001010011110011000010101000010011010010100000011010001011101111110000110001100011010001001101111110,
128'b0000110000010010011001100110001001001001011001111010001000110101110010001110110100101100100100011001001100100111110001111110010,
128'b1011100111001111010100111110111100111110010001011111011100111001010101000110111100000011001010101110010011001000101101000110111,
128'b0110001110010000110111011111101100010010000110011001101010001000011110111000010101110000110010001101101100101100000011011101111,
128'b1100010101000100011110101111101100001000010101101111101010100110000100010110000000000011011000000110001101010100100000110000000,
128'b0010000010111111101100011111010110110100111100111010111101101111000001011100010010101011000011011000000001011100010011101000111,
128'b0011111011100000000101100000011011010010101101111101000110000100111010110110010101001011110111010110110111000001111111010001010,
128'b1011111001111101000101011110001000011001111011000001010101100000111011011010111001000000011101000111110111110000011010110110100,
128'b1000011011010000001011110011100011000101010101110110100100100001000000010101000010001101111010101110100111000001000100111001001,
128'b0000000100100111011100001010111100010111111101111000110001100111010101010000101011000100011010111111111111101010011010100010000,
128'b0100011011001101000110101100111011001011110010000000010110011101110001100001100110000110000110000000010110111111111000111111100,
128'b0000111111000100001011111110101011110100001110001111011010010110100100000000110110000001001110110101111010101011011110100110010,
128'b1101101001110111111100101100010101100101010000000011001111011100010101011100010110000110010111000000110011110100101100010100010,
128'b0110000000100111111001111001100001011001000001011010011100000111000100001011101010111011110100001000101110000111001100100100100,
128'b0000010101000100011010010010011110000111101111101100000000000110100011011111000011100101100000111100000000100000100111001011101,
128'b1010101100111110001110011101111010011111110110110100110000001110110000111101100011101010111100101010010000111011101110001100100,
128'b0101110101011011011111001101101000001101100111101111001110101010000110101101110101101111000100100101010011010000111111001110111,
128'b0100001001110101001000100100101011111011110001011110000101101111111100100001111010101100001110010000110010100111111101011010010,
128'b1101011010001111111000000101001110000000100011101111010000111101001111011111111101011010001000001011110011001110011101111101100,
128'b1110100010001011010110110010111101010100100000010010011000100100000111011001000110010111101101011111110000101010110100100111001,
128'b1011011111011110110010001010011000000000001111101011011111001010100011111001010101110011110111010101101000100110000100110000000,
128'b1000000110011110010001100011111110011101110000010100010101001111100000011001101001010001000111101100010001110101101010010100001,
128'b0000101111100011000010101000101000000001101000100000111111100011100000010000100001101110110010111100001101010111110001001000101,
128'b0100100110110110011100111011010011100011111001101101111111011001110011110110101101111111110010011110110010010110111000000001001,
128'b1001100010000100001100010010110010001100010100101010110111001011101001010111100000110100010011110011011101111100011101011011010,
128'b0101101100001110010111011000101101001100100000111100000110111001110100011001100011011101101111010100110111101001001101111111010,
128'b0001101110110111000000010011011101010011110101000001110001000000101101111001111001001010110001101001000011100110001101010011010,
128'b0101010010010010011011111001011001001110001110111000000100001100011000100011010101000110111111100001101011100111001100000011001,
128'b1001000010000001111010010001010101001001001100110010011111011111010100001001111100100001101111100110001011111010010010101111000,
128'b0001100111011011010000110110010011110101110100000000111110011000001110011100100110001101010000000101110101110011010011010111000,
128'b0100011101011011100010001001101000101100011001100100000111000100011000111001000011110001010010010101001101111110111101010000100,
128'b1101101010000101010100110000011101111000011011000000101000111100011101001100010010000110110111101001001101000001000100100111000,
128'b1010101111111100001100001100000011001111000000000100001010111100000010111111010101111010110110110111011001001011100001010011101,
128'b0000010111000100111011011011101100011100010011111011110000001100011100101011001110011110101010100001100010010001111111100011000,
128'b1101101010111001111101001100010101010110101011101001110101010100000010011010110010111010111011100100100000110010001111011101111,
128'b0001110110010010101000110001100001110100111000001000001100010011010101101111111110110011100001111000010010000010011010100010000,
128'b1111100110011101101001000011100011101001100111110100001100010101110001010010111000000100001010010100011000110000111100010010100,
128'b1100010001011111010010010101111010101100010110001011001010101001001111001111100010110101001101000110101110110010010110100011101,
128'b0011110001000110011110011111110000010001100010010011001110100011100110111101111011111111011001110001001111000010000001001111001,
128'b0011111101101111000011100111000101011101101100010001011101010101110011110101011110111011000001110110111111010000100110001001000,
128'b1110011100001000111011001111110010111101011110000001110101101100001010001101001011111000110101111011001010010101000111010100111,
128'b0001111001111000010001000011001100101110010110110111101110101001111010010011001001111110000000111001100110110111111100111101110,
128'b0011000111100110110010101100100110101110011011000100011010001110000101011001001010111101110111110001000111000011011111101011100,
128'b0001010101000101001000011101011011011001101100001100111101111010010010100011001111010001001110100111100100010011010111010011010,
128'b1100001000010100100110111001011010010101110010100001010010111001001000001011100101010011110000100101100111101100000000101101111,
128'b1100000101000110001110110010010111100001010011110100010100011010011101101000100100000001111010100000010101101000101100011101010,
128'b1101110110001100010111011111010000100011001100010101010111101110101100100011011011110000100000110001001101100111100100100111000,
128'b0010001000100001000110100000001100010010001001000111101001000111110110110110011100010010101111101010000110000110111001011110001,
128'b1010011101011001110100001001110110100111101111110111100111001100100110110010111100111000010101111110100011111011111000010010001,
128'b0100110000100110111011010000110010110011100010010011111011101110000110111110000101101101000100111010010010000101110110011010000,
128'b0011100010001010100000110110101111011101000010100111110011110010110011111110110001000011001011100011001110100111011110111111110,
128'b1100101110110000010101000011010110000100100111100111110001011111010110100101000010001011011011100000100000111100101010101010101,
128'b1111111011101010110001101000101101011100010111001111010101011010100001100001100111111110110110110101111100000110010001011111011,
128'b0101101010101110001111111101100001000101001010110110011001100100010111010001011001101100000100011011010111111100011011011001010,
128'b1000100110111101011101010001101101000101100100011111010111011000001000000011001111111000010110011011001011001011011001010111001,
128'b0010011101100001110101100001110100110110010001110001110000001111010110101001111111010010010011000010110110001011101000110110110,
128'b0111010001101010001100110110010000010110101100010101111001101000000110001010011100001100010001000110110110010011100001011110110,
128'b1110101100000001101001000101011111001000100000010010011010100100000011110110000101101011101100101111101111011001110100000111110,
128'b1000100011000100100111100000110101010000110111011111111110111001011001000110000110000110110100110110000011111001110110101110000,
128'b1011011001100111111001011010010010010011011010101101111110111111110101011111101110111110111000101011111011011101010000000010010,
128'b0111001100001001001101001011100010101000111100100000011001001101011001010111100010101010001100101111100000010111011011101111000,
128'b1111110000111111010110000000001011100010110101000100101000100111111100011001101001010000011110011011000100000011101001011111111,
128'b1111000100111001010001101100010101111000011110110010001111110110010111000011100010110010110111011100011111001111010011010110000,
128'b0011011111101100010100100111010001110111101000001101110010011000101111100000000010111101110100000110111100101111011101101001111,
128'b1100011101111011111000010111100100001001000110011011101000011010110000100011010101001000001000101001000111001000010101110001101,
128'b0110111010110101111101000001100101001110100011000000100001111100001110001101110101100011001000101000011011101101000010110001100,
128'b0100011010000001110010010101001011010110100001110101000100000000001101101111100001100111111010101011000100011111111000011101110,
128'b1110100000111101001010011110011110011111101101111010010010100100100100001000101100111100111110011011001111011010001110001110110,
128'b1011100000011101001111001011011110110011111000101111111111010111111011111101000011110100001011001111111011000101001011101010000,
128'b0101101110010011101101001011010001011011001101101111001001101100101000010111001110001111111110001111011000101101100001010011100,
128'b1010001010111011110010111101000101100000011111000100011001111001011000000100110101100001110011101000000001111101110000010110000,
128'b0001001111110101000100011100101100111100100011100000011110110000110011011001011111111011000111100011011100011001101011101010001,
128'b1010011110001010101001010001001101011110110001101110110101111110101111111000010000100011001001000110111010111101111100110010010,
128'b1111010100010001101101010000000000111101010111011001100010001000111110010001111111000101101101011101010011100100101000110101000,
128'b0100011011110000110001010010010110101101001100100010111011010101001011111100111011100101000000001000100110111101001011101001010,
128'b0101011010111100011100100000001111100001111001111011110011110111100010010110010011010111001111101001010010011110001011100011111,
128'b0101110111110101001110101011000011011110101011101110101110001111110100011001001110000011011010010010110110100011110001110101110,
128'b0001101010101100111110101111101111101001111111001101001010110100011101110101011001101100100101010110111011110010101000011011010,
128'b0100011101100110010000000011010011100100011001100010000010101011101110001110000100001000010111110100001100110111001001100101001,
128'b1010110110000010011000110011001000010100101110010111101100101101001001011100010111111101010010111001101000001101011000101000101,
128'b0011101101000001111101001000101101001110111110101100111000000001100010110100010011000110111000111011101101100101111000010001100,
128'b0110001110000111111110111000011000100000011011110000000101101100110011111110110010001101000111010101010010101011100101011100010,
128'b1001010110100111100101111010111110100101000010101010110001111101000000011101010101110100011111100110011010101011110010100100000,
128'b0101100011010011000111010010101111110100100011100000110101010010100010010110010011111111110110101001001000110100010100111001011,
128'b1100001101101110010001111100110011011100000100011001111110100000000000000011001100110110001010100100111000111100110110000111000,
128'b0001110001111110000011010001111101111000101111111110000110101101110001011100001010100100111111011101100100110011010010110011111,
128'b1011111000111110000011000110101101010110110111001011000110110110100000001101010110011110110010100000010110001001000101001000110,
128'b1010100001110110001110010111111000000000001101000000101101000110100011101010001110101111101111111101001110000101000000000011000,
128'b1101100101000110011000110111101101110010101011010011000101100001101110000000011101001101100001000101010001111001001000110101000,
128'b0011101111110011001100000001001101101011100001110000001010100111100011010111010100011111001000010011011100011010111001001000000,
128'b1110010001011010110110100111000111111001100100110111001101010011010001101010101110000010110101100011111011011000100110111111001,
128'b1001011010100000110011100111101101110101110011001100111110110111111011001001111101010000001001001000100000010000011111010100111,
128'b1001000000000011111111110011110101000100000001100111011111000111111010101001001110011010110011000101110001111101110101011001100,
128'b1101011111100100001101010100011001010001011111010111011010111001110001011110001100011011101111110000001111010101111001100101001,
128'b0101110000001101101011101110101101110000000100010111101000011000100111000110001001010100111010010001000011110110000111100101001,
128'b1010000111000001001001011001100001100010001101010010101110111100100011011110100110010101010001000010101111000110110010100000101,
128'b1110101010001010111111010000111010000110010101011011001010101100000100111011101001111100100110001010110111011000100000110110110,
128'b1111101101100100011100101100000111100101110010010001100110110010011001010101101001011110000110100000011001111010111101110000100,
128'b0010111111011011010100110100111110011110011111001101010011110001000101010010001010110010010001111101000100000011000011010101010,
128'b1011011110110011001111100001111110011100110010101010101111100011001011111100011111110000110001000100101001110001010000101010100,
128'b0001000100110001010000101010111001001000011100001110010010010000110000110100010101111010100001001111010001111000110011111011110,
128'b0110111001000010101100110101111011010001111001111001000010100111010111001101010000110111000000010010111011110101001010010000101,
128'b0111010000100100101101001101000100111110000111001101101011100010001101111100001000110101100111100111111001010000000010010010101,
128'b1110010011001100111001110111110011100011111110101100010011110011100011011110010000001011101010111100011110111111101111001011001,
128'b0101100010101101010011010110010001101000000110111101111100001110100000011100110110001111000110110000101101101001110110001000010,
128'b0010100100111001111111001111000101010101011000010111000010110111000101111100110110011101000101110001010010000111100001010101000,
128'b0110110110000000010101110111111000110101100111111101001100000111111101000101110001110110010011101000100011000100111101000101010,
128'b1110000101101011000000110111001011001011010011100000011000010100101010101110110011001101011101101000100000000101111101000000011,
128'b1111101100000111101110000010000111001110100000111101100010000010100111010011011110111101000010100110011000110011100011110010100,
128'b1000110111010010101001111101110101111111111111111001011111111101001000010010100010101011011001010011000100101101101110000000000,
128'b1111010111010010101011010111011011101100001001000010000011000011110100111100001100000000010001001100000110110000010010111001100,
128'b1010000101001101000000010101100110111001111010010111100001010101011011110110010100110001110110111001101001101001010010111101011,
128'b1111011111000110001101100101110100010100010001000011100111110100101000111100000000000100001111010100100101000000111011100101111,
128'b1010001000100100101100100100100000010010001001100001000100001111111011110011011011001010010100010111010100100000100001011111011,
128'b0011000010101100000111111010010011110000110000110101100000100100010001110001101001011110000001000111001001100000010101111101000,
128'b0110110111011000001011010010000110110100101110101001001101010100110100101000011001011101011000110000010000111110000111000111010,
128'b1100111101010100101111000000111100111011111110110101011011110011011001001001110101010110001101100110010101001101001000111111001,
128'b0100001101010001101000001000101110000100001111101010100000100110110110000001011101101010100111011111001111001010101000101100010,
128'b0101100001001001000011000111101110000100010111000100111101111111000010011111010101010011111111011011010011111110010000001010000,
128'b0010010100011111011011000110001100010111111110101110111010000111101110011000010100110101011011010001000010111111101000101010000,
128'b0111010011101011110010010001010111000011100001011011111000100101100111010100000110000000001111110010001001011010111110110001111,
128'b0100101100001010000001100001011110001100111111100001011001111100100000000011011001111101011101101010010101000101010101011110001,
128'b1010001110110111000010001111110111000010101110011010101111101011110101001000011100000010000100100000000010101111100111101100001,
128'b1011010001110010100001001110010010111101111111110110010011000101110001100110111100111111100110001111101101111011011011100101111,
128'b0011101011110001101011110010100011010111111110110010010011101101010000010110000000000100000010010011100111001100011001101101101,
128'b1001111001101111100110100101100100001101000010010110110000110111101011010011101000101111111101011110111000000110111110011101111,
128'b0101010100000100011110111111000100111011000101011011010001011001111000011111001110101010000110001100111001011101011001010011101,
128'b1011011011010100011011111101110110111101101110100100100100000111101010011100011010000001111000111000111101111101001011101001001,
128'b1010011100001111011011001110110110101110101001110001010011100001110010000001101111100011111110111000011111001010001010011001011,
128'b0000100000010101000100001110110010110000000110110100001101110111111101011101000110111011010001000111000101010110010000111100010,
128'b0010011111000100100111001100100001101111101010011001001000000000111110111001110100000111100111010010011001000000011101001110111,
128'b0000100100011100010001101101010010000100001001100001101110011000011000101100100101110111011111001010111000011000101000110001001,
128'b1100001011010000011010100111110100001101010101110000000110100000110010010101101010100000100100011001100001100111010100000010101,
128'b0110011000001000000111010001111011001001100111110100110110100111000011011110001100111100010001001000010100100111011101111000011,
128'b1011010011000101000111000011001000111001000010101000010000101100010111110101110110010100100000011111100001100000101101001110111,
128'b0100111111001011100010001001011001110100110010111110011011010100010101111011000011001010111001011101000100100000110101001111010,
128'b0100000101111110110001010001100101110101100011000111010010111001001000101000011111111100010000001111101111001010100010000110010,
128'b1001001001000011011000010010111100100111011000101111110111111001010011010001000000001101101000000000011100101101111100000110100,
128'b0110001111100010010001101100101010000000100111011001001110000100100010010101111011111111000101111111100011001011010100001111001,
};
