module target_word(input [6:0] index, output [24:0] word);

localparam [24:0] wordlist [0:99] = {
25'b0011100010100110000001100, //match
25'b1000110100011000010001011, //lemur
25'b0010010010100011010001111, //purse
25'b0111001000100011010000010, //curio
25'b0101100100001001001110010, //steel
25'b1100001011010110111000111, //holly
25'b1001110111010001011010011, //twixt
25'b1100000011101000000000110, //gaudy
25'b0101100000110000111001011, //loyal
25'b0101101000101010010000011, //devil
25'b1100010011100110100000011, //ditty
25'b1001110010010001011010011, //twist
25'b0101010010010001000100101, //frisk
25'b1001110001001001010101110, //overt
25'b0011100010100111010000001, //butch
25'b0101001101101000101100101, //flunk
25'b0010010010000000000100000, //abase
25'b0010000010010001011010011, //twice
25'b0101000010000000101100001, //black
25'b1100000100000100100000011, //dicey
25'b1011100000100010111000001, //borax
25'b0111101100101000011100010, //chump
25'b1000100100011110010001011, //leper
25'b1011001110100011000100000, //arrow
25'b1000100100000110001101110, //odder
25'b1100010011100110000000001, //batty
25'b0001100000001000011100000, //ahead
25'b1001110100000010010010001, //rebut
25'b1001110010010000111000111, //hoist
25'b0011101111011001010000111, //humph
25'b1100001100010000101110010, //slimy
25'b0001100100010110000100000, //abled
25'b1000110100011100101100101, //flour
25'b1100001011110000000000110, //gayly
25'b0010010101000001010010010, //suave
25'b1000100100010100000010011, //taker
25'b0101000010011100110010010, //smock
25'b0010000011011100000100000, //abode
25'b1000100100101110100000101, //fixer
25'b1100000100001100000000010, //cagey
25'b1100010001010000000000111, //hairy
25'b1001010100000100100000101, //ficus
25'b0010010100000010110001000, //imbue
25'b0110100000011000111010110, //woman
25'b0111010001100110110101000, //intro
25'b0011110011010000000000101, //faith
25'b0010010010001000010000110, //geese
25'b1001101011000000010000011, //dealt
25'b1100010011000000010001100, //meaty
25'b1001100000001000011110110, //wheat
25'b0011110011011100111010010, //sooth
25'b1001100010010001010100100, //evict
25'b1001010010110000000100000, //abyss
25'b1011000100010101001000000, //askew
25'b1000100100101010010000101, //fever
25'b0010010010010111010001111, //pulse
25'b0010000010010001000110011, //trice
25'b0101001101101000101101111, //plunk
25'b1001101101001001010100100, //event
25'b0011001101010000111000110, //going
25'b1100001011010111010010010, //sully
25'b0101000010001000101100101, //fleck
25'b0010010001011100001010010, //score
25'b0001101101101000111001100, //mound
25'b1001110100011100000100000, //about
25'b1100001101011100011101111, //phony
25'b1011001110000110100010110, //widow
25'b1100010011001010010001011, //lefty
25'b1000101110000010000001011, //labor
25'b1001100100001001000100110, //greet
25'b0010010001011010010000110, //genre
25'b1000100100000010110000000, //amber
25'b0011100010100110010010001, //retch
25'b1100001110101010000010010, //savoy
25'b0011100010011010000010001, //ranch
25'b1100001011010110111000110, //golly
25'b0101001101000000101100001, //blank
25'b0110101110010110010001100, //melon
25'b0111101000010111010010011, //tulip
25'b0011100010010000011110110, //which
25'b0010010010011101000101111, //prose
25'b0111101100101001000100010, //crump
25'b0011100110101000111000011, //dough
25'b1100000101001010100001001, //jiffy
25'b0010010001001000011110110, //where
25'b0011100110101000000001011, //laugh
25'b0010001100011100110100110, //gnome
25'b0000101100010000101100010, //climb
25'b1001100101011100101100000, //aloft
25'b0101101000000000101100101, //flail
25'b0010001111011100101110010, //slope
25'b0101100000000100010000101, //fecal
25'b0010010101000001000100010, //crave
25'b0101100000100010100010101, //viral
25'b1100001011101100111001011, //lowly
25'b0010001000100010010000100, //eerie
25'b1000101110000111000100000, //ardor
25'b1000100100001001001110010, //steer
25'b1100001101011101000101000, //irony
25'b0010001101011100101100000 //alone
};

assign word = wordlist[index];

endmodule
