module word_db (input [24:0] word, input clk, input rst, output wire in_db);

//Bloom filter storing 1000 words in 4096 bits with 4 hash functions
localparam [11:0] hash_params [0:3] [0:4] = {
{12'h01a5, 12'h06b3, 12'h0e6c, 12'h0dd0, 12'h0c0f},
{12'h04fc, 12'h0f69, 12'h0874, 12'h05ce, 12'h09ae},
{12'h036e, 12'h0c84, 12'h0c0a, 12'h060a, 12'h028f},
{12'h0663, 12'h0c61, 12'h0dfe, 12'h0724, 12'h0cfb}
};

(* ramstyle = "block" *) localparam bloom_filter [0:4095] = {
64'b110011111110000011111110001111000101100000000011101110110101111,
64'b011110110111110011011110111000001111101111010101010111000110111,
64'b111011000010011111101110111110101111011110001011000111110000101,
64'b101100111110101011100111011111100111101101110001111010100101111,
64'b111110011011011000111111111111001100111010010110101110110100101,
64'b000100011111101101111110010100100111101101100010000111101111111,
64'b011110100101111111011101100000011001100011110001011110111110011,
64'b010101001101110010111011111101110111101100011111000010110111001,
64'b011111100001110100110000011101010011001110100010101111100010110,
64'b011111101011111011100111001111111110011010100111001101111010110,
64'b111101100010111100110001101111001110110101001110001111001100011,
64'b011011100111101111001001111001101110111101110111111000110011011,
64'b011010011011000011100000111111101011011100010001101001110100011,
64'b111010011101111101011001100111001001001111001010111000110010110,
64'b011111101010100010111111010111100111010110111101101001100110100,
64'b100011010101110101111011100111101111011111011001110010110101110,
64'b110110101101011010110110110011001010011111010111111001001111111,
64'b011010110011111110111011101111010100111100100101111100101011110,
64'b000111011011101010001001001011100011010001101011101111101101100,
64'b111111011111001110101110011111000110101011111001000010110101101,
64'b111111111110100010110100110000011011101111111011111101100000100,
64'b010110001100111110001001011100101011111010010000111111000000110,
64'b010101110110110111000111010101100010110010111110011111101011100,
64'b101100111001101110110111111000001011001001111011011110111011111,
64'b011101101111000001011101111001010111010101011011111011111010111,
64'b011111100001111110010001101111110001100010101111111111100011110,
64'b111001111000111111111011100110011010111011011010000111101111101,
64'b111001000110101101100010010110000111111110011111111111011101101,
64'b100111111110101010101110111010111101111110100111111001111111101,
64'b111111001100101111100111111101000111011011000001111011111101100,
64'b000100101001111110011111111011111101110100011111001110101010011,
64'b111111111101110001110110101111100011111100100001100011101110010,
64'b111110101111101111111111010101110101010010101111101011010001111,
64'b011111111101001111100100001011010011100110001110100011101010111,
64'b011010110111111111001101111001110110110111011111001010101110111,
64'b001001110011011110101010111111100100010110111110111100111110011,
64'b010011101111011000111010110101001100100110101000110001111000111,
64'b100101111111111111001111111001101010001111101100011100100111010,
64'b110011011000111110111001111011111001001111011000111101111101110,
64'b111110101001101110010110100010001111111010000001111111110011101,
64'b111111100100111010100110111111011110111011101110000111100111101,
64'b010010100010111110111010111000100101001111100101100100110010110,
64'b111011110111011111101111101111101110001111110011101000100111111,
64'b010111111000001111010000111111100011011001111010100110110010010,
64'b101001110001111110101101011011001100011011101011000010100110100,
64'b101101111011010011010011100100010011101111011111101110111010011,
64'b011110110111101111101110110010010111010001000101101111101101011,
64'b010110100111101111011110011011010011011011100111101111111111100,
64'b011001001011100111100001111011011111001011110001101110011010000,
64'b011100111111100110101111110001100110001100001110101011101111011,
64'b111010111101111110000110111000011110111101100100011011111101101,
64'b100111101011111110111110100111011011100101111010111101100111111,
64'b001000011101111100110010101111011101111101111100101000101011101,
64'b111110111011011111111111011110101011011001101000011110111101010,
64'b011111111110101100001101001111101101011001111100000100101101111,
64'b111001000111101101010111011011111111011010101100111001000101111,
64'b100111000100110110010010001111011001001110100100010111100010111,
64'b110111110010000010110010110010110101110111001101101111111001111,
64'b101010110100110010111010101110001110111111111100011111100111001,
64'b011111111010001001110111011011100110011011111001100101100000101,
64'b010000001011111011100010111101111010111011111010110101011011110,
64'b100100101111111101000100111001001110101101101100110010110001111,
64'b001111001111111001111001111111001111110110001110010010101111111,
64'b100111101100101111110010111110110001101101000000111001111000100
};

wire [11:0] hash_table [0:4];

wire [11:0] hash;

reg [0:3] in_db_i;

reg [1:0] i;

genvar j;
generate
for (j = 0; j < 5; j = j + 1) begin : which_letter
assign hash_table[j] = hash_params[i][j] * word[5*j + 4:5*j];
end
endgenerate
assign hash = hash_table[0] + hash_table[1] + hash_table[2] + hash_table[3] + hash_table[4];

always @(posedge clk or posedge rst) begin
    if (rst) begin
        i <= 0;
        in_db_i <= 4'b0;
    end else begin
        i <= i+1;
    end
end
        
assign in_db_i[i] = bloom_filter[hash[i]];

assign in_db = &in_db_i;

endmodule
